module and_gate(input g_input, e_input, output o);
	assign o = g_input & e_input;
endmodule
